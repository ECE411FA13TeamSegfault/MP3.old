--
-- VHDL Architecture ece411.NOT1.untitled
--
-- Created:
--          by - schen79.ews (linux-a2.ews.illinois.edu)
--          at - 13:12:41 09/20/13
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY NOT1 IS
   PORT( 
      A : IN     std_logic;
      F : OUT    std_logic
   );

-- Declarations

END NOT1 ;

--
ARCHITECTURE untitled OF NOT1 IS
BEGIN
	PROCESS(A)
		VARIABLE NOTInternal : std_logic;
		BEGIN
			NOTInternal := NOT A;
			F <= NOTInternal after DELAY_LOGIC2;
		END PROCESS;
END ARCHITECTURE untitled;

